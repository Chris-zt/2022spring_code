module shifter
	#(parameter N = 8,
	  RST_VALUE = {N{1'b0}})
	  


endmodule