module counter 
	#(parameter N = 8,
	RST_VALUE = {N{1'b1}})
	(input clk, rst, pe, ce,
	input [N-1:0]
	
	);
	
endmodule