module nmux2 (
	ports
);
	
endmodule