module register (
	input rst, clk, en,
	input [31:0] d,
	output [31:0] q
);
	
	
endmodule