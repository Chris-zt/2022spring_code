module Adder (
	ports
);
	
endmodule