module Adder (
	input [3:0] Ln, [15:0] Out,
	output add
);
	wire
	
endmodule